`ifndef __SQUAT_HEADER__

`define __SQUAT_HEADER__

`define CHANNEL_NUM 16

`endif