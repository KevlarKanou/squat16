`ifndef __SQUART_HEADER__

`define __SQUART_HEADER__

`define CHANNEL_NUM 16

`endif