`ifndef __SQUAT_HEADER__

`define __SQUAT_HEADER__

`define PORT_NUM 16

`endif