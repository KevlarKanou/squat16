`ifndef __SQUAT_HEADER__

`define __SQUAT_HEADER__

`define PORT_NUM        16

`define UNI_VPI_WIDTH   8
`define UNI_VCI_WIDTH   16

`define NNI_VPI_WIDTH   12
`define NNI_VCI_WIDTH   16

`define ForwardLoc      43:28
`define NNIVPILoc       27:16
`define NNIVCILoc       15:0

`endif